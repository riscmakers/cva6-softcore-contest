
`define ARIANE_DATA_WIDTH 64

// Instantiate protocl checker
// `define PROTOCOL_CHECKER

// write-back cache
// `define WB_DCACHE

// write-through cache
//`define WT_DCACHE

// RISC Makers data cache
`define RISCMAKERS_DCACHE

// debug probe
//`define LAUTERBACH_DEBUG_PROBE

// to use DDR connecting to Zynq PS  
`define PS7_DDR


